`timescale 1ns/1ps

module FPCVT_tb;

  logic [11:0] D;
  logic        S;
  logic [2:0]  E;
  logic [3:0]  F;

  FPCVT dut (
    .D(D),
    .S(S),
    .E(E),
    .F(F)
  );
    
    initial begin
    automatic logic [11:0] patterns [0:34] = '{
        12'b0000_0000_0000,
        12'b1111_1111_1111,
        12'b0000_0000_0001,
        12'b1000_0000_0000,
        12'b0101_0101_0101,
        12'b0111_1111_1111,
        12'b0111_1111_0001,
        12'b0000_0000_1000,
        12'b0100_1110_0101,
        12'b0010_1011_0011,
        12'b1010_1010_1010,
        12'b1100_0000_0000,
        12'b0010_1100_1000,
        12'b0111_1110_1111,
        12'b0011_1100_0000,
        12'b1110_0001_1010,
        12'b0001_0010_1111,
        12'b0000_0001_0001, 
        12'b0000_0010_0010, 
        12'b0000_0100_0100,
        12'b0000_1000_1000, 
        12'b0010_0000_0001, 
        12'b0011_0000_0011, 
        12'b0100_0000_1111, 
        12'b0100_1001_0000, 
        12'b0110_0110_0110, 
        12'b0110_1110_1110, 
        12'b1001_0001_0001, 
        12'b1011_1000_1000, 
        12'b1101_0101_0101, 
        12'b1110_1110_0000, 
        12'b1111_0000_1111, 
        12'b1111_1000_0001, 
        12'b0111_0001_1110,
        12'b0011_1110_0000
    };

        foreach (patterns[i]) begin
            D = patterns[i];
            #10; 
            $display("[%0t] D = %b | S = %b | E = %d | F = %b",
                     $time, D, S, E, F);
        end
    $finish;
    end
endmodule
